LIBRARY IEEE;
--USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CLK_1HZ IS
	PORT (
		MCLK : IN BIT;
		CLKOUT : OUT BIT
	);
END CLK_1HZ;

ARCHITECTURE Behavioral OF CLK_1HZ IS
	SIGNAL COUNTER : INTEGER RANGE 0 TO 24_999_999 := 0;
	SIGNAL C1HZ : BIT;
BEGIN
	PROCESS (MCLK)
	BEGIN
		IF MCLK = '1' AND MCLK'EVENT THEN
			IF COUNTER = 24_999_999 THEN
				COUNTER <= 0;
				C1HZ <= NOT C1HZ;
			ELSE COUNTER <= COUNTER + 1;
			END IF;
		ELSE NULL;
		END IF;
	END PROCESS;

	CLKOUT <= C1HZ;
END Behavioral;