--Stephanie Denisse Benitez Cabrera
--Práctica 4
--Segundo componente (decoder)

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity BCDto4Display is
    Port ( BCD_in : in STD_LOGIC_VECTOR (3 downto 0);
           LED_out : out STD_LOGIC_VECTOR (6 downto 0));
end  BCDto4Display;

architecture arch of  BCDto4Display is
begin
process(BCD_in)
    begin
        case BCD_in is
        when "0000" => LED_out <= "0000001"; -- "0"     
        when "0001" => LED_out <= "1001111"; -- "1" 
        when "0010" => LED_out <= "0010010"; -- "2" 
        when "0011" => LED_out <= "0000110"; -- "3" 
        when "0100" => LED_out <= "1001100"; -- "4" 
        when "0101" => LED_out <= "0100100"; -- "5" 
        when "0110" => LED_out <= "0100000"; -- "6" 
        when "0111" => LED_out <= "0001111"; -- "7" 
        when "1000" => LED_out <= "0000000"; -- "8"     
        when "1001" => LED_out <= "0000100"; -- "9" 
        when others => null;
        end case;
    end process;
        end arch;